// system verilog implmentation of a memory controller
// uses cache.sv and ram.sv