// system verilog implmentation of a cache