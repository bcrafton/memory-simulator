// system verilog implementation of a memory controller
// uses cache.sv and ram.sv